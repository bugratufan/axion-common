--------------------------------------------------------------------------------
-- Axion Common Library
-- 
-- Shared VHDL modules and utilities for Axion FPGA projects.
-- 
-- Copyright (c) 2024 Bugra Tufan
-- MIT License
--------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

library work;
use work.axion_common_pkg.all;

package axion_common is
    -- This package provides access to all axion_common components
    -- See individual source files for component declarations
end package axion_common;
